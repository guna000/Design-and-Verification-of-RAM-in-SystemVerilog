parameter DATA_WIDTH = 8;
parameter ADDR_BUS_WIDTH = 6 ;
parameter MAX_MEM_LOC = (2**ADDR_BUS_WIDTH)-1;
parameter MAX_DATA_VAL = (2**(DATA_WIDTH-1))-1;